module ucmp1(a, b : sup, equ)
	equ = a*b + /a*/b
  sup = a*/b
end module
